interface fa();
  logic in_a,in_b,in_cin;
  logic sum,carry;
endinterface
