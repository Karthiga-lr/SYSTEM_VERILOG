interface inti();
logic a;
logic b;
logic cin;
logic s;
logic cout;

endinterface
