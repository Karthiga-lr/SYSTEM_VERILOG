interface intf;
  logic clk;
  logic rst;
  logic d;
  logic [3:0] count;
endinterface
