module int_example;
  int i;
  initial begin 
    i = 123496;
    $display("int: %0d", i);
  end
endmodule
