// To _Do
