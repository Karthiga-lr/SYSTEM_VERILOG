///TO-DO
