// TO D
