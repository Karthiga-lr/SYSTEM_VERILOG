//TO - DO
