module assoc_array_find;
