module AND_gate(input a,input b, input clk, output y);
  assign y = a && b;
endmodule
