// to -do
